LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
ENTITY ALU2 IS
PORT (Clock :in std_logic; --input clock signal
		A,B :in unsigned (7 downto 0); -- 8 bit inputs from latches A and B
		student_id : in unsigned (3 downto 0); --4 bit student id from fsm
		OP: in unsigned (15 downto 0); --16 bit selector for Operation from Decorder
		Neg: out std_logic; --is the result negative? se -ve bit output
		R1 : out unsigned(3 downto 0); --lower 4 bits of 8 bit result output
		R2 : out unsigned(3 downto 0)); --higher 4 bits of 8 bi result output
end ALU2;
architecture calculation of ALU2 is --temporary signal declrations
signal Reg1, Reg2, Result : unsigned(7 downto 0):=(others=> '0');
signal Reg4 : unsigned (0 to 7);
begin 
Reg1<=A; --temporarily store A in Reg1 local vairable
Reg2<=B; --temporarily store B in Reg2 local variable 
process (Clock,OP)
begin	
	if (rising_edge(Clock)) THEN --Do the calculation @positive edge of clock
	case OP is
		WHEN "0000000000000001" =>
			--Decrement by 9
			Result<=(Reg2)-9;
		WHEN "0000000000000010" => --Swap the lower and upper 4 bits of B
			Result (3 downto 0)<= B(7 downto 4);
			Result (7 downto 4)<= B(3 downto 0);
		WHEN "0000000000000100"=> --Shift A to left by 2 bits
			Result<=Reg1 sll 2;
		WHEN "0000000000001000"=>--NANDing A and B
			Result<= Reg1 NAND Reg2;
		WHEN "0000000000010000"=>--Find greater value of A and B and produce result
			if (Reg1>Reg2) then
				Result<=Reg1;
				end if;
			if (Reg2>Reg1) then
				Result<=Reg2;
				end if;
		WHEN "0000000000100000" => --Invert even bits of B
			Result<= NOT B;
		WHEN "0000000001000000"=>--Produce null on the output
			Result<= null;
		WHEN "0000000010000000"=>--Replace the upper four bits of B by upper four bits of A
			Result (7 downto 4)<= Reg1 (7 downto 4) ;
			Result (3 downto 0)<= Reg2(3 downto 0);
		WHEN "0000000100000000" =>--Show A on the output
			Result<= Reg1;
		WHEN OTHERS =>
			--Dont care, do nothing
end case;
end if;
end process;
R1 <= Result (3 downto 0);
R2 <= Result (7 downto 4);
end calculation;